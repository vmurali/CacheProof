typedef Bit#(TLog#(n)) Bitt#(type n);
typedef Bit#(TLog#(TAdd#(n, 1))) NumElems#(type n);
